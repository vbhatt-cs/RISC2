library ieee;
use ieee.std_logic_1164.all;
package mem_package is
type ram_t is array (0 to 255) of std_logic_vector(15 downto 0);
constant INST_INIT : ram_t := (
0 => "1000000000011101",
1 => "0100100110000101",
2 => "0001110000111101",
3 => "0100110110000101",
4 => "0110000000000011",
5 => "0001000010000000",
6 => "0010000001011000",
7 => "0010011011011000",
8 => "0001011011000000",
9 => "0000100010100001",
10 => "0000000000000000",
11 => "0010110110110010",
12 => "1100110101111010",
13 => "0101100101010110",
29 => "0001011011000001",
30 => "0001110110010111",
31 => "0001001001011111",
32 => "0001001001001110",
33 => "0101000110000100",
34 => "0100000110000000",
35 => "1100101001001100",
36 => "0000000010010000",
37 => "0000011100100010",
38 => "0001001001111111",
39 => "0001111111111100",
47 => "0001110000000010",
48 => "0111000000010100",
49 => "0001011011111111",
50 => "0101011110000101",
51 => "0100111110000100",
others => (others => '0'));

constant DATA_INIT : ram_t := (
20 => x"0001",
21 => x"000F",
--22 => x"000C",
23 => x"FFFF",
24 => x"0045",
--25 => x"FFBB",
--26 => x"0044",
others => (others => '0'));
end package mem_package;